module my_or (output y, input a, b);
	or or1(y, a, b);
endmodule 