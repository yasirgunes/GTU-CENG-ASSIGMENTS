module myAdd(input A, B, output C);

assign C = A & B;






endmodule
