// my_and

module my_and(output result, input a, b);
	and and1 (result, a, b);
endmodule