module small_m(A, B, Y);
input A;
input B;
output Y;

assign Y = A & B;


endmodule
