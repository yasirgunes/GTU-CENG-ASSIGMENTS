// my_or 

module my_or (output result, input a, b);
	or or1 (result, a, b);
endmodule 