module extend_to_32(output [31:0] result, input a);

and and1(result[0], a, 1);
and and2(result[1], a, 1);
and and3(result[2], a, 1);
and and4(result[3], a, 1);
and and5(result[4], a, 1);
and and6(result[5], a, 1);
and and7(result[6], a, 1);
and and8(result[7], a, 1);
and and9(result[8], a, 1);
and and10(result[9], a, 1);
and and11(result[10], a, 1);
and and12(result[11], a, 1);
and and13(result[12], a, 1);
and and14(result[13], a, 1);
and and15(result[14], a, 1);
and and16(result[15], a, 1);
and and17(result[16], a, 1);
and and18(result[17], a, 1);
and and19(result[18], a, 1);
and and20(result[19], a, 1);
and and21(result[20], a, 1);
and and22(result[21], a, 1);
and and23(result[22], a, 1);
and and24(result[23], a, 1);
and and25(result[24], a, 1);
and and26(result[25], a, 1);
and and27(result[26], a, 1);
and and28(result[27], a, 1);
and and29(result[28], a, 1);
and and30(result[29], a, 1);
and and31(result[30], a, 1);
and and32(result[31], a, 1);

endmodule
