module my_and (output y, input a, b);
	and and1(y, a, b);
endmodule 