module and_31bit(
    output [30:0] result,
    input [30:0] A,
    input [30:0] B
);

and and1(result[0], A[0], B[0]);
and and2(result[1], A[1], B[1]);
and and3(result[2], A[2], B[2]);
and and4(result[3], A[3], B[3]);
and and5(result[4], A[4], B[4]);
and and6(result[5], A[5], B[5]);
and and7(result[6], A[6], B[6]);
and and8(result[7], A[7], B[7]);
and and9(result[8], A[8], B[8]);
and and10(result[9], A[9], B[9]);
and and11(result[10], A[10], B[10]);
and and12(result[11], A[11], B[11]);
and and13(result[12], A[12], B[12]);
and and14(result[13], A[13], B[13]);
and and15(result[14], A[14], B[14]);
and and16(result[15], A[15], B[15]);
and and17(result[16], A[16], B[16]);
and and18(result[17], A[17], B[17]);
and and19(result[18], A[18], B[18]);
and and20(result[19], A[19], B[19]);
and and21(result[20], A[20], B[20]);
and and22(result[21], A[21], B[21]);
and and23(result[22], A[22], B[22]);
and and24(result[23], A[23], B[23]);
and and25(result[24], A[24], B[24]);
and and26(result[25], A[25], B[25]);
and and27(result[26], A[26], B[26]);
and and28(result[27], A[27], B[27]);
and and29(result[28], A[28], B[28]);
and and30(result[29], A[29], B[29]);
and and31(result[30], A[30], B[30]);


endmodule
