module deneme (input a, b, c, output [31:0] d);
assign d[0] = a&b;

endmodule
